//Deassert the wrreq signal in the same clock cycle when the full signal is asserted.
//Deassert the rdreq signal in the same clock cycle when the empty signal is asserted.
//
module Chn_fifo_Control
(
  input clk,
  input reset_n,
  input rst_all_fifo,
  input [15:0] chn1_Dataout,
  input chn1_Dataout_en,
  input [15:0] chn2_Dataout,
  input chn2_Dataout_en,
  output reg [15:0] out_to_usb_ext_fifo_din,
  output reg out_to_usb_ext_fifo_en
);
//chn1
reg chn1_fifo_empty;
reg chn1_fifo_full;
reg chn1_fifo_rdreq;
reg [15:0] chn1_out_to_usb_fifo;
reg [10:0] chn1_fifo_usedw;
sync_fifo chn1_fifo
(
	aclr(~reset_n | rst_all_fifo),
	clock(clk),
	data(chn1_Dataout),
	wrreq(chn1_Dataout_en & (!chn2_fifo_full)),
	empty(chn1_fifo_empty),
	full(chn1_fifo_full),
	rdreq(chn1_fifo_rdreq),  
	q(chn1_out_to_usb_fifo),
	usedw(chn1_fifo_usedw)
);
//chn2
reg chn2_fifo_empty;
reg chn2_fifo_full;
reg chn2_fifo_rdreq;
reg [15:0] chn2_out_to_usb_fifo;
reg [10:0] chn2_fifo_usedw;
sync_fifo chn2_fifo
(
	aclr(~reset_n | rst_all_fifo),
	clock(clk),
	data(chn2_Dataout),
	wrreq(chn2_Dataout_en & (!chn2_fifo_full)),
	empty(chn2_fifo_empty),
	full(chn2_fifo_full),
	rdreq(chn2_fifo_rdreq),  
	q(chn2_out_to_usb_fifo),
	usedw(chn2_fifo_usedw)
);
always @ (posedge clk , negedge reset_n) begin
  if(!reset_n) begin
    chn1_fifo_empty = 1'b0;
    chn1_fifo_full = 1'b0;
    chn1_rdreq = 1'b0;
    [15:0] chn1_out_to_usb_fifo = 16'h0;
    [10:0] chn1_usedw = 11'b000_0000_0000;
    chn2_fifo_empty = 1'b0;
    chn2_fifo_full = 1'b0;
    chn2_rdreq = 1'b0;
    [15:0] chn2_out_to_usb_fifo = 16'h0000;
    [10:0] chn2_usedw = 11'b000_0000_0000;
  end
end 
//ѡ���ȡ��һ��FIFO�����ݣ�ÿ�ζ���һ��FIFO��Ͷ�����һ��FIFO
parameter Chn1_fifo_selected = 1'b0;
          Chn2_fifo_selected = 1'b1;
reg Select_State;
reg fifo_rdreq;
//reg fifo_full;
//reg fifo_empty;
reg [15:0] fifo_buffer;
reg [10:0] fifo_usedw;
always @ (posedge clk , negedge reset_n) begin
  if (~reset_n) begin
    Select_State <= Chn1_fifo_selected;
    fifo_rdreq <= 1'b0;
    //fifo_full <= 1'b0;
    //fifo_empty <= 1'b0;
    fifo_buffer <= 16'h0;
    fifo_usedw <= 11'b0;
  end
  else begin
    case (Select_State)
      Chn1_fifo_selected:begin
        chn1_fifo_rdreq <= fifo_rdreq;
        //fifo_full <= chn1_fifo_full;
        //fifo_empty <= chn1_fifo_empty;
        fifo_buffer <= chn1_out_to_usb_fifo;
        fifo_usedw <= chn1_fifo_used;
      end
      Chn2_fifo_selected:begin 
        chn2_fifo_rdreq <= fifo_rdreq;
        //fifo_full <= chn2_fifo_full;
        //-fifo_empty <= chn2_fifo_empty;
        fifo_buffer <= chn2_out_to_usb_fifo;
        fifo_usedw <= chn2_fifo_usedw;
      end 
  end
//fifo��ȡ����
parameter fifo_read_num = 10'd1023;//ÿ�ζ�fifo��һ��������������һ��fifoʱ��֤����һ��fifo��Ҫװ��
reg [9:0] fifo_read_cnt;//
parameter [2:0] IDLE = 3'd0;
                CHECK = 3'd1;
                WAIT = 3'd2;
                READ = 3'd3;
                WAIT_DONE = 3'd4;
                DONE = 3'd5;
reg [2:0] State;
always @ (posedge clk , negedge reset_n) begin
  if(~reset_n) begin
    fifo_rdreq <=  1'b0;
    fifo_usedw <= 11'd0;
    fifo_buffer <= 16'h0;
  end
  else begin
    case(State)
      IDLE:
        fifo_raed_cnt <= 10'b0;
        State <= CHECK;
      CHECK:begin
        if(fifo_usedw > fifo_read_num) begin

      end
  end


end


endmodule
